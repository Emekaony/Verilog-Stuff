/*
this is the test bench for the half adder
*/

`include "/Users/shadon./Developer/verilog_stuff/src/half_adder.v"

module half_adder_tb;
    reg a, b;

    // to declare output use wire
    wire sum, carry;

    half_adder add1(a, b, sum, carry);

    initial begin
        // dump the changes in of the code
        // vcd means value changed dump
        $dumpfile("half_adder.vcd");
        $dumpvars(0, half_adder_tb);

        a=0; b=0;
        #1
        a=0; b=1;
        #1
        a=1; b=0;
        #1
        a=1; b=1;
    end

endmodule